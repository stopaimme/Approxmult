module approxmult_16bits (
    input wire [15:0] INA,INB,
    output wire [31:0] result
);
    wire [19:0]sig;
    wire [15:0]a,b;
    reg [15:0] p[15:0];
    sub s(.a({4'b0000,INA}),.diff({4,b0000,INB}),.s(sig),.co());
    assign a = sig[19]?INB:INA;
    assign b = sig[19]?INA:INB;
    integer i,j;
    always@(*)begin
        for(i = 0; i<=15; i = i + 1)
            for(j = 0; j <= 15; j = j + 1)
                p[i][j] = a[j] & b[i];
    end   

    
//----------------Partial product generation----------------
    wire [2:0] s1[35:0];
    half_add h1(p[0][8],p[1][7],s1[0][0],s1[0][1]);

    ap_comp ap1(p[0][9],p[1][8],p[2][7],p[3][6],s1[1][0],s1[1][1]);

    ap_comp ap2(p[0][10],p[1][9],p[2][8],p[3][7],s1[2][0],s1[2][1]);
    half_add h2(p[4][6],p[5][5],s1[3][0],s1[3][1]);

    ap_comp ap3(p[0][11],p[1][10],p[2][9],p[3][8],s1[4][0],s1[4][1]);
    ap_comp ap4(p[4][7],p[5][6],p[6][5],p[7][4],s1[5][0],s1[5][1]); 

    ap_comp ap5(p[0][12],p[1][11],p[2][10],p[3][9],s1[6][0],s1[6][1]);
    ap_comp ap6(p[4][8],p[5][7],p[6][6],p[7][5],s1[7][0],s1[7][1]);
    half_add h3(p[8][4],p[9][3],s1[8][0],s1[8][1]);

    ap_comp ap7(p[0][13],p[1][12],p[2][11],p[3][10],s1[9][0],s1[9][1]);
    ap_comp ap8(p[4][9],p[5][8],p[6][7],p[7][6],s1[10][0],s1[10][1]);
    ap_comp ap9(p[8][5],p[9][4],p[10][3],p[11][2],s1[11][0],s1[11][1]);

    ap_comp ap10(p[0][14],p[1][13],p[2][12],p[3][11],s1[12][0],s1[12][1]);
    ap_comp ap11(p[4][10],p[5][9],p[6][8],p[7][7],s1[13][0],s1[13][1]);
    ap_comp ap12(p[8][6],p[9][5],p[10][4],p[11][3],s1[14][0],s1[14][1]);
    half_add h4(p[12][2],p[13][1],s1[15][0],s1[15][1]);

    ap_comp ap13(p[0][15],p[1][14],p[2][13],p[3][12],s1[16][0],s1[16][1]);
    ap_comp ap14(p[4][11],p[5][10],p[6][9],p[7][8],s1[17][0],s1[17][1]);
    ap_comp ap15(p[8][7],p[9][6],p[10][5],p[11][4],s1[18][0],s1[18][1]);
    ap_comp ap16(p[12][3],p[13][2],p[14][1],p[15][0],s1[19][0],s1[19][1]);

    ap_comp ap17(p[1][15],p[2][14],p[3][13],p[4][12],s1[20][0],s1[20][1]);
    ap_comp ap18(p[5][11],p[6][10],p[7][9],p[8][8],s1[21][0],s1[21][1]);
    ap_comp ap19(p[9][7],p[10][6],p[11][5],p[12][4],s1[22][0],s1[22][1]);
    half_add h5(p[13][3],p[14][2],s1[23][0],s1[23][1]);

    ap_comp ap20(p[2][15],p[3][14],p[4][13],p[5][12],s1[24][0],s1[24][1]);
    ap_comp ap21(p[6][11],p[7][10],p[8][9],p[9][8],s1[25][0],s1[25][1]);
    ap_comp ap22(p[10][7],p[11][6],p[12][5],p[13][4],s1[26][0],s1[26][1]);

    ap_comp ap23(p[3][15],p[4][14],p[5][13],p[6][12],s1[27][0],s1[27][1]);
    ap_comp ap24(p[7][11],p[8][10],p[9][9],p[10][8],s1[28][0],s1[28][1]);
    half_add h6(p[11][7],p[12][6],s1[29][0],s1[29][1]);

    ap_comp ap25(p[4][15],p[5][14],p[6][13],p[7][12],s1[30][0],s1[30][1]);
    ap_comp ap26(p[8][11],p[9][10],p[10][9],p[11][8],s1[31][0],s1[31][1]);

    ap_comp ap27(p[5][15],p[6][14],p[7][13],p[8][12],s1[32][0],s1[32][1]);
    half_add h7(p[9][11],p[10][10],s1[33][0],s1[33][1]);
    

    ap_comp ap28(p[6][15],p[7][14],p[8][13],p[9][12],s1[34][0],s1[34][1]);

    half_add h8(p[7][15],p[8][14],s1[35][0],s1[35][1]);

//----------------Partial product reduction1----------------
    wire [2:0] s2[38:0];
    ap_comp ap29(p[2][6],p[3][5],p[4][4],s1[0][0],s2[0][0],s2[0][1]);
    ap_comp ap30(p[5][3],p[6][2],p[7][1],p[8][0],s2[1][0],s2[1][1]);

    ap_comp ap31(p[4][5],p[5][4],s1[1][0],s1[0][1],s2[2][0],s2[2][1]);
    ap_comp ap32(p[6][3],p[7][2],p[8][1],p[9][0],s2[3][0],s2[3][1]);

    ap_comp ap33(p[6][4],s1[2][0],s1[3][0],s1[1][1],s2[4][0],s2[4][1]);
    ap_comp ap34(p[7][3],p[8][2],p[9][1],p[10][0],s2[5][0],s2[5][1]);

    ap_comp ap35(s1[4][0],s1[5][0],s1[2][1],s1[3][1],s2[6][0],s2[6][1]);
    ap_comp ap36(p[8][3],p[9][2],p[10][1],p[11][0],s2[7][0],s2[7][1]);

    ap_comp ap37(s1[6][0],s1[7][0],s1[4][1],s1[5][1],s2[8][0],s2[8][1]);
    ap_comp ap38(p[10][2],p[11][1],p[12][0],s1[8][0],s2[9][0],s2[9][1]);

    ap_comp ap39(s1[9][0],s1[10][0],s1[6][1],s1[7][1],s2[10][0],s2[10][1]);
    ap_comp ap40(s1[11][0],s1[8][1],p[12][1],p[13][0],s2[11][0],s2[11][1]);

    ap_comp ap41(s1[12][0],s1[13][0],s1[9][1],s1[10][1],s2[12][0],s2[12][1]);
    ap_comp ap42(s1[14][0],s1[15][0],s1[11][1],p[14][0],s2[13][0],s2[13][1]);

    ap_comp ap43(s1[16][0],s1[17][0],s1[12][1],s1[13][1],s2[14][0],s2[14][1]);
    ap_comp ap44(s1[18][0],s1[19][0],s1[14][1],s1[15][1],s2[15][0],s2[15][1]);

    ap_comp ap45(s1[20][0],s1[21][0],p[15][1],s1[17][1],s2[16][0],s2[16][1]);
    ap_comp ap46(s1[22][0],s1[23][0],s1[18][1],s1[19][1],s2[17][0],s2[17][1]);

    ap_comp ap47(s1[24][0],s1[25][0],p[14][3],s1[22][1],s2[18][0],s2[18][1]);
    ap_comp ap48(s1[26][0],s1[21][1],p[15][2],s1[23][1],s2[19][0],s2[19][1]);

    ap_comp ap49(s1[27][0],s1[28][0],p[13][5],s1[25][1],s2[20][0],s2[20][1]);
    ap_comp ap50(s1[29][0],p[14][4],p[15][3],s1[26][1],s2[21][0],s2[21][1]);

    ap_comp ap51(s1[30][0],p[12][7],p[13][6],s1[28][1],s2[22][0],s2[22][1]);
    ap_comp ap52(s1[31][0],p[14][5],p[15][4],s1[29][1],s2[23][0],s2[23][1]);

    ap_comp ap53(s1[32][0],p[11][9],p[12][8],p[13][7],s2[24][0],s2[24][1]);
    ap_comp ap54(s1[33][0],p[14][6],p[15][5],s1[31][1],s2[25][0],s2[25][1]);

    ap_comp ap55(s1[34][0],p[10][11],p[11][10],p[12][9],s2[26][0],s2[26][1]);
    ap_comp ap56(p[13][8],p[14][7],p[15][6],s1[33][1],s2[27][0],s2[27][1]);

    ap_comp ap57(s1[35][0],p[9][13],p[10][12],p[11][11],s2[28][0],s2[28][1]);
    ap_comp ap58(p[12][10],p[13][9],p[14][8],p[15][7],s2[29][0],s2[29][1]);

    ac_comp ac1(p[8][15],p[9][14],p[10][13],p[11][12],1'b0,s2[30][0],s2[30][1],s2[30][2]);
    ac_comp ac2(p[12][11],p[13][10],p[14][9],p[15][8],1'b0,s2[31][0],s2[31][1],s2[31][2]);

    ac_comp ac3(p[9][15],p[10][14],p[11][13],p[12][12],s2[30][2],s2[32][0],s2[32][1],s2[32][2]);
    ac_comp ac4(p[13][11],p[14][10],p[15][9],1'b0,s2[31][2],s2[33][0],s2[33][1],s2[33][2]);
    
    ac_comp ac5(p[10][15],p[11][14],p[12][13],p[13][12],s2[32][2],s2[34][0],s2[34][1],s2[34][2]);
    add a1(p[14][11],p[15][10],s2[33][2],s2[35][0],s2[35][1]);

    ac_comp ac6(p[11][15],p[12][14],p[13][13],p[14][12],s2[34][2],s2[36][0],s2[36][1],s2[36][2]);

    add a2(p[12][15],p[13][14],s2[36][2],s2[37][0],s2[37][1]);

    Err_detect E1(p[10][12],p[11][11],p[14][8],p[15][7],s2[38][0]);

//----------------Partial product reduction2------------------
    wire [2:0] s3[21:0];

    half_add h9(s2[0][0],s2[1][0],s3[0][0],s3[0][1]);

    ap_comp ap59(s2[0][1],s2[1][1],s2[2][0],s2[3][0],s3[1][0],s3[1][1]);

    ap_comp ap60(s2[2][1],s3[3][1],s3[4][0],s3[5][0],s3[2][0],s3[2][1]);

    ap_comp ap61(s2[4][1],s2[5][1],s2[6][0],s2[7][0],s3[3][0],s3[3][1]);

    ap_comp ap62(s2[6][1],s2[7][1],s2[8][0],s2[9][0],s3[4][0],s3[4][1]);

    ap_comp ap63(s2[8][1],s2[9][1],s2[10][0],s2[11][0],s3[5][0],s3[5][1]);

    ap_comp ap64(s2[10][1],s2[11][1],s2[12][0],s2[13][0],s3[6][0],s3[6][1]);

    ap_comp ap65(s2[12][1],s2[13][1],s2[14][0],s2[15][0],s3[7][0],s3[7][1]);

    ap_comp ap66(s2[14][1],s2[15][1],s2[16][0],s2[17][0],s3[8][0],s3[8][1]);

    ap_comp ap67(s2[16][1],s2[17][1],s2[18][0],s2[19][0],s3[9][0],s3[9][1]);

    ap_comp ap68(s2[18][1],s2[19][1],s2[20][0],s2[21][0],s3[10][0],s3[10][1]);

    ap_comp ap69(s2[20][1],s2[21][1],s2[22][0],s2[23][0],s3[11][0],s3[11][1]);

    ap_comp ap70(s2[22][1],s2[23][1],s2[24][0],s2[25][0],s3[12][0],s3[12][1]);

    ap_comp ap71(s2[24][1],s2[25][1],s2[26][0],s2[27][0],s3[13][0],s3[13][1]);

    ap_comp ap72(s2[26][1],s2[27][1],s2[28][0],s2[29][0],s3[14][0],s3[14][1]);

    ac_comp ac7(1'b0,1'b0,s2[30][0],s2[31][0],s2[38][0],s3[15][0],s3[15][1],s3[15][2]);

    ac_comp ac8(s2[30][1],s2[31][1],s2[32][0],s2[33][0],s3[15][2],s3[16][0],s3[16][1],s3[16][2]);

    ac_comp ac9(s2[32][1],s2[33][1],s2[34][0],s2[35][0],s3[16][2],s3[17][0],s3[17][1],s3[17][2]);

    ac_comp ac10(s2[34][1],s2[35][1],s2[36][0],p[15][11],s3[17][2],s3[18][0],s3[18][1],s3[18][2]);

    ac_comp ac11(s2[36][1],s2[37][0],p[14][13],p[15][12],s3[18][2],s3[19][0],s3[19][1],s3[19][2]);

    ac_comp ac12(s2[37][1],p[13][15],p[14][14],p[15][13],s3[19][2],s3[20][0],s3[20][1],s3[20][2]);

    add a3(p[14][15],p[15][14],s3[20][2],s3[21][0],s3[21][1]);


//----------------Carry propagation adder------------------

    wire [1:0] s4[21:0];

    half_add h10(s3[0][1],s3[1][0],s4[0][0],s4[0][1]);

    add a4(s3[1][1],s3[2][0],s4[0][1],s4[1][0],s4[1][1]);

    add a5(s3[2][1],s3[3][0],s4[1][1],s4[2][0],s4[2][1]);

    add a6(s3[3][1],s3[4][0],s4[2][1],s4[3][0],s4[3][1]);

    add a7(s3[4][1],s3[5][0],s4[3][1],s4[4][0],s4[4][1]);

    add a8(s3[5][1],s3[6][0],s4[4][1],s4[5][0],s4[5][1]);

    add a9(s3[6][1],s3[7][0],s4[5][1],s4[6][0],s4[6][1]);

    add a10(s3[7][1],s3[8][0],s4[6][1],s4[7][0],s4[7][1]);

    add a11(s3[8][1],s3[9][0],s4[7][1],s4[8][0],s4[8][1]);

    add a12(s3[9][1],s3[10][0],s4[8][1],s4[9][0],s4[9][1]);

    add a13(s3[10][1],s3[11][0],s4[9][1],s4[10][0],s4[10][1]);

    add a14(s3[11][1],s3[12][0],s4[10][1],s4[11][0],s4[11][1]);

    add a15(s3[12][1],s3[13][0],s4[11][1],s4[12][0],s4[12][1]);

    add a16(s3[13][1],s3[14][0],s4[12][1],s4[13][0],s4[13][1]);

    add a17(s3[14][1],s3[15][0],s4[13][1],s4[14][0],s4[14][1]);

    add a18(s3[15][1],s3[16][0],s4[14][1],s4[15][0],s4[15][1]);

    add a19(s3[16][1],s3[17][0],s4[15][1],s4[16][0],s4[16][1]);

    add a20(s3[17][1],s3[18][0],s4[16][1],s4[17][0],s4[17][1]);

    add a21(s3[18][1],s3[19][0],s4[17][1],s4[18][0],s4[18][1]);

    add a22(s3[19][1],s3[20][0],s4[18][1],s4[19][0],s4[19][1]);

    add a23(s3[20][1],s3[21][0],s4[19][1],s4[20][0],s4[20][1]);

    add a24(s3[21][1],p[15][15],s4[20][1],s4[21][0],s4[21][1]);






    
    assign result[0] = 1'b0;
    assign result[1] = 1'b0;
    assign result[2] = 1'b0;
    assign result[3] = 1'b0;
    assign result[4] = 1'b0;
    assign result[5] = 1'b0;
    assign result[6] = 1'b0;
    assign result[7] = 1'b0;
    assign result[8] = s3[3][0];
    assign result[9] = s4[0][0];
    assign result[10] = s4[1][0];
    assign result[11] = s4[2][0];
    assign result[12] = s4[3][0];
    assign result[13] = s4[4][0];
    assign result[14] = s4[5][0];
    assign result[15] = s4[6][0];
    assign result[16] = s4[7][0];
    assign result[17] = s4[8][0];
    assign result[18] = s4[9][0];
    assign result[19] = s4[10][0];
    assign result[20] = s4[11][0];
    assign result[21] = s4[12][0];
    assign result[22] = s4[13][0];
    assign result[23] = s4[14][0];
    assign result[24] = s4[15][0];
    assign result[25] = s4[16][0];
    assign result[26] = s4[17][0];
    assign result[27] = s4[18][0];
    assign result[28] = s4[19][0];
    assign result[29] = s4[20][0];
    assign result[30] = s4[21][0];
    assign result[31] = s4[21][1];

endmodule